.title SRAM_6T_CORE_16x8_MC_TB
.include /home/majh/OpenYield/sim/20260124_224745_mc_6t/tmp_mc.spice
.param U=0
.DC U -0.71 0.71 0.001
.SAMPLING useExpr=true
.options samples numsamples=1
.PRINT DC FORMAT=NOINDEX {U} V(V1) V(V2)
.subckt SRAM_6T_CELL_DISCONNECT VDD VSS BL BLB WL
MPGL BL WL QD VSS NMOS_VTG l=5e-08 w=1.35e-07
MPGR BLB WL QBD VSS NMOS_VTG l=5e-08 w=1.35e-07
MPDL QD QB VSS VSS NMOS_VTG l=5e-08 w=9e-08
MPDR QBD Q VSS VSS NMOS_VTG l=5e-08 w=9e-08
MPUL QD QB VDD VDD PMOS_VTG l=5e-08 w=9e-08
MPUR QBD Q VDD VDD PMOS_VTG l=5e-08 w=9e-08
.ends SRAM_6T_CELL_DISCONNECT
VVDD VDD VSS 1.0V
VVSS VSS 0 0V
XSRAM_6T_CELL_DISCONNECT VDD VSS BL BLB WL SRAM_6T_CELL_DISCONNECT
VWL_gnd WL VSS 0V
EV1 V1 VSS VOL='U+sqrt(2)*V(XSRAM_6T_CELL_DISCONNECT:QBD)'
EV2 V2 VSS VOL='-U+sqrt(2)*V(XSRAM_6T_CELL_DISCONNECT:QD)'
EQ XSRAM_6T_CELL_DISCONNECT:Q VSS  VOL='1/sqrt(2)*U+1/sqrt(2)*V(V1)'
EQB XSRAM_6T_CELL_DISCONNECT:QB VSS  VOL='-1/sqrt(2)*U+1/sqrt(2)*V(V2)'
EVD VD VSS VOL='ABS(V(V1)-V(V2))'
.options TEMP = 27C
.options TNOM = 27C
.ic V(BL)=1.0V V(BLB)=1.0V
.meas DC MAXVD MAX V(VD)
.meas DC HOLD_SNM PARAM='1/sqrt(2)*MAXVD'
.end
