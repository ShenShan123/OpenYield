.title SRAM_6T_CORE_16x8_MC_TB
.include /home/majh/OpenYield/sim/20260124_204333_mc_6t/tmp_mc.spice
.TRAN 1.0000e-11 5.0000e-09
.OPTIONS OUTPUT INITIAL_INTERVAL=1.0000e-11
.SAMPLING useExpr=true
.options samples numsamples=1
.PRINT TRAN FORMAT=NOINDEX V(CLK) V(CLK_BUF) V(CLK_BAR) V(CSB) V(CS_BAR) V(CS) V(WEB) V(WE_BAR) V(WE) V(GATED_CLK_BUF) V(GATED_CLK_BAR) V(WL_EN) V(RWL)
.PRINT TRAN FORMAT=NOINDEX V(A0) V(A_DFF0) V(A1) V(A_DFF1) V(A2) V(A_DFF2) V(A3) V(A_DFF3) V(RBL) V(RBL_DELAY) V(RBL_DELAY_BAR) V(W_EN) V(PRE)
.PRINT TRAN FORMAT=NOINDEX V(S_EN) V(WL15) V(BL7) V(BLB7) V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_15_7:Q) V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_15_7:QB) 
.PRINT TRAN V(SA_Q7) V(SA_QB7)V(OUT)
.subckt SRAM_6T_CORE_16x8 VDD VSS BL0 BL1 BL2 BL3 BL4 BL5 BL6 BL7 BLB0 BLB1 BLB2 BLB3 BLB4 BLB5 BLB6 BLB7 WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15
.subckt SRAM_6T_CELL VDD VSS BL BLB WL
MPGL BL WL Q VSS NMOS_VTG l=5e-08 w=1.35e-07
MPGR BLB WL QB VSS NMOS_VTG l=5e-08 w=1.35e-07
MPDL Q QB VSS VSS NMOS_VTG l=5e-08 w=9e-08
MPDR QB Q VSS VSS NMOS_VTG l=5e-08 w=9e-08
MPUL Q QB VDD VDD PMOS_VTG l=5e-08 w=9e-08
MPUR QB Q VDD VDD PMOS_VTG l=5e-08 w=9e-08
.ends SRAM_6T_CELL
XSRAM_6T_CELL_0_0 VDD VSS BL0 BLB0 WL0 SRAM_6T_CELL
XSRAM_6T_CELL_0_1 VDD VSS BL1 BLB1 WL0 SRAM_6T_CELL
XSRAM_6T_CELL_0_2 VDD VSS BL2 BLB2 WL0 SRAM_6T_CELL
XSRAM_6T_CELL_0_3 VDD VSS BL3 BLB3 WL0 SRAM_6T_CELL
XSRAM_6T_CELL_0_4 VDD VSS BL4 BLB4 WL0 SRAM_6T_CELL
XSRAM_6T_CELL_0_5 VDD VSS BL5 BLB5 WL0 SRAM_6T_CELL
XSRAM_6T_CELL_0_6 VDD VSS BL6 BLB6 WL0 SRAM_6T_CELL
XSRAM_6T_CELL_0_7 VDD VSS BL7 BLB7 WL0 SRAM_6T_CELL
XSRAM_6T_CELL_1_0 VDD VSS BL0 BLB0 WL1 SRAM_6T_CELL
XSRAM_6T_CELL_1_1 VDD VSS BL1 BLB1 WL1 SRAM_6T_CELL
XSRAM_6T_CELL_1_2 VDD VSS BL2 BLB2 WL1 SRAM_6T_CELL
XSRAM_6T_CELL_1_3 VDD VSS BL3 BLB3 WL1 SRAM_6T_CELL
XSRAM_6T_CELL_1_4 VDD VSS BL4 BLB4 WL1 SRAM_6T_CELL
XSRAM_6T_CELL_1_5 VDD VSS BL5 BLB5 WL1 SRAM_6T_CELL
XSRAM_6T_CELL_1_6 VDD VSS BL6 BLB6 WL1 SRAM_6T_CELL
XSRAM_6T_CELL_1_7 VDD VSS BL7 BLB7 WL1 SRAM_6T_CELL
XSRAM_6T_CELL_2_0 VDD VSS BL0 BLB0 WL2 SRAM_6T_CELL
XSRAM_6T_CELL_2_1 VDD VSS BL1 BLB1 WL2 SRAM_6T_CELL
XSRAM_6T_CELL_2_2 VDD VSS BL2 BLB2 WL2 SRAM_6T_CELL
XSRAM_6T_CELL_2_3 VDD VSS BL3 BLB3 WL2 SRAM_6T_CELL
XSRAM_6T_CELL_2_4 VDD VSS BL4 BLB4 WL2 SRAM_6T_CELL
XSRAM_6T_CELL_2_5 VDD VSS BL5 BLB5 WL2 SRAM_6T_CELL
XSRAM_6T_CELL_2_6 VDD VSS BL6 BLB6 WL2 SRAM_6T_CELL
XSRAM_6T_CELL_2_7 VDD VSS BL7 BLB7 WL2 SRAM_6T_CELL
XSRAM_6T_CELL_3_0 VDD VSS BL0 BLB0 WL3 SRAM_6T_CELL
XSRAM_6T_CELL_3_1 VDD VSS BL1 BLB1 WL3 SRAM_6T_CELL
XSRAM_6T_CELL_3_2 VDD VSS BL2 BLB2 WL3 SRAM_6T_CELL
XSRAM_6T_CELL_3_3 VDD VSS BL3 BLB3 WL3 SRAM_6T_CELL
XSRAM_6T_CELL_3_4 VDD VSS BL4 BLB4 WL3 SRAM_6T_CELL
XSRAM_6T_CELL_3_5 VDD VSS BL5 BLB5 WL3 SRAM_6T_CELL
XSRAM_6T_CELL_3_6 VDD VSS BL6 BLB6 WL3 SRAM_6T_CELL
XSRAM_6T_CELL_3_7 VDD VSS BL7 BLB7 WL3 SRAM_6T_CELL
XSRAM_6T_CELL_4_0 VDD VSS BL0 BLB0 WL4 SRAM_6T_CELL
XSRAM_6T_CELL_4_1 VDD VSS BL1 BLB1 WL4 SRAM_6T_CELL
XSRAM_6T_CELL_4_2 VDD VSS BL2 BLB2 WL4 SRAM_6T_CELL
XSRAM_6T_CELL_4_3 VDD VSS BL3 BLB3 WL4 SRAM_6T_CELL
XSRAM_6T_CELL_4_4 VDD VSS BL4 BLB4 WL4 SRAM_6T_CELL
XSRAM_6T_CELL_4_5 VDD VSS BL5 BLB5 WL4 SRAM_6T_CELL
XSRAM_6T_CELL_4_6 VDD VSS BL6 BLB6 WL4 SRAM_6T_CELL
XSRAM_6T_CELL_4_7 VDD VSS BL7 BLB7 WL4 SRAM_6T_CELL
XSRAM_6T_CELL_5_0 VDD VSS BL0 BLB0 WL5 SRAM_6T_CELL
XSRAM_6T_CELL_5_1 VDD VSS BL1 BLB1 WL5 SRAM_6T_CELL
XSRAM_6T_CELL_5_2 VDD VSS BL2 BLB2 WL5 SRAM_6T_CELL
XSRAM_6T_CELL_5_3 VDD VSS BL3 BLB3 WL5 SRAM_6T_CELL
XSRAM_6T_CELL_5_4 VDD VSS BL4 BLB4 WL5 SRAM_6T_CELL
XSRAM_6T_CELL_5_5 VDD VSS BL5 BLB5 WL5 SRAM_6T_CELL
XSRAM_6T_CELL_5_6 VDD VSS BL6 BLB6 WL5 SRAM_6T_CELL
XSRAM_6T_CELL_5_7 VDD VSS BL7 BLB7 WL5 SRAM_6T_CELL
XSRAM_6T_CELL_6_0 VDD VSS BL0 BLB0 WL6 SRAM_6T_CELL
XSRAM_6T_CELL_6_1 VDD VSS BL1 BLB1 WL6 SRAM_6T_CELL
XSRAM_6T_CELL_6_2 VDD VSS BL2 BLB2 WL6 SRAM_6T_CELL
XSRAM_6T_CELL_6_3 VDD VSS BL3 BLB3 WL6 SRAM_6T_CELL
XSRAM_6T_CELL_6_4 VDD VSS BL4 BLB4 WL6 SRAM_6T_CELL
XSRAM_6T_CELL_6_5 VDD VSS BL5 BLB5 WL6 SRAM_6T_CELL
XSRAM_6T_CELL_6_6 VDD VSS BL6 BLB6 WL6 SRAM_6T_CELL
XSRAM_6T_CELL_6_7 VDD VSS BL7 BLB7 WL6 SRAM_6T_CELL
XSRAM_6T_CELL_7_0 VDD VSS BL0 BLB0 WL7 SRAM_6T_CELL
XSRAM_6T_CELL_7_1 VDD VSS BL1 BLB1 WL7 SRAM_6T_CELL
XSRAM_6T_CELL_7_2 VDD VSS BL2 BLB2 WL7 SRAM_6T_CELL
XSRAM_6T_CELL_7_3 VDD VSS BL3 BLB3 WL7 SRAM_6T_CELL
XSRAM_6T_CELL_7_4 VDD VSS BL4 BLB4 WL7 SRAM_6T_CELL
XSRAM_6T_CELL_7_5 VDD VSS BL5 BLB5 WL7 SRAM_6T_CELL
XSRAM_6T_CELL_7_6 VDD VSS BL6 BLB6 WL7 SRAM_6T_CELL
XSRAM_6T_CELL_7_7 VDD VSS BL7 BLB7 WL7 SRAM_6T_CELL
XSRAM_6T_CELL_8_0 VDD VSS BL0 BLB0 WL8 SRAM_6T_CELL
XSRAM_6T_CELL_8_1 VDD VSS BL1 BLB1 WL8 SRAM_6T_CELL
XSRAM_6T_CELL_8_2 VDD VSS BL2 BLB2 WL8 SRAM_6T_CELL
XSRAM_6T_CELL_8_3 VDD VSS BL3 BLB3 WL8 SRAM_6T_CELL
XSRAM_6T_CELL_8_4 VDD VSS BL4 BLB4 WL8 SRAM_6T_CELL
XSRAM_6T_CELL_8_5 VDD VSS BL5 BLB5 WL8 SRAM_6T_CELL
XSRAM_6T_CELL_8_6 VDD VSS BL6 BLB6 WL8 SRAM_6T_CELL
XSRAM_6T_CELL_8_7 VDD VSS BL7 BLB7 WL8 SRAM_6T_CELL
XSRAM_6T_CELL_9_0 VDD VSS BL0 BLB0 WL9 SRAM_6T_CELL
XSRAM_6T_CELL_9_1 VDD VSS BL1 BLB1 WL9 SRAM_6T_CELL
XSRAM_6T_CELL_9_2 VDD VSS BL2 BLB2 WL9 SRAM_6T_CELL
XSRAM_6T_CELL_9_3 VDD VSS BL3 BLB3 WL9 SRAM_6T_CELL
XSRAM_6T_CELL_9_4 VDD VSS BL4 BLB4 WL9 SRAM_6T_CELL
XSRAM_6T_CELL_9_5 VDD VSS BL5 BLB5 WL9 SRAM_6T_CELL
XSRAM_6T_CELL_9_6 VDD VSS BL6 BLB6 WL9 SRAM_6T_CELL
XSRAM_6T_CELL_9_7 VDD VSS BL7 BLB7 WL9 SRAM_6T_CELL
XSRAM_6T_CELL_10_0 VDD VSS BL0 BLB0 WL10 SRAM_6T_CELL
XSRAM_6T_CELL_10_1 VDD VSS BL1 BLB1 WL10 SRAM_6T_CELL
XSRAM_6T_CELL_10_2 VDD VSS BL2 BLB2 WL10 SRAM_6T_CELL
XSRAM_6T_CELL_10_3 VDD VSS BL3 BLB3 WL10 SRAM_6T_CELL
XSRAM_6T_CELL_10_4 VDD VSS BL4 BLB4 WL10 SRAM_6T_CELL
XSRAM_6T_CELL_10_5 VDD VSS BL5 BLB5 WL10 SRAM_6T_CELL
XSRAM_6T_CELL_10_6 VDD VSS BL6 BLB6 WL10 SRAM_6T_CELL
XSRAM_6T_CELL_10_7 VDD VSS BL7 BLB7 WL10 SRAM_6T_CELL
XSRAM_6T_CELL_11_0 VDD VSS BL0 BLB0 WL11 SRAM_6T_CELL
XSRAM_6T_CELL_11_1 VDD VSS BL1 BLB1 WL11 SRAM_6T_CELL
XSRAM_6T_CELL_11_2 VDD VSS BL2 BLB2 WL11 SRAM_6T_CELL
XSRAM_6T_CELL_11_3 VDD VSS BL3 BLB3 WL11 SRAM_6T_CELL
XSRAM_6T_CELL_11_4 VDD VSS BL4 BLB4 WL11 SRAM_6T_CELL
XSRAM_6T_CELL_11_5 VDD VSS BL5 BLB5 WL11 SRAM_6T_CELL
XSRAM_6T_CELL_11_6 VDD VSS BL6 BLB6 WL11 SRAM_6T_CELL
XSRAM_6T_CELL_11_7 VDD VSS BL7 BLB7 WL11 SRAM_6T_CELL
XSRAM_6T_CELL_12_0 VDD VSS BL0 BLB0 WL12 SRAM_6T_CELL
XSRAM_6T_CELL_12_1 VDD VSS BL1 BLB1 WL12 SRAM_6T_CELL
XSRAM_6T_CELL_12_2 VDD VSS BL2 BLB2 WL12 SRAM_6T_CELL
XSRAM_6T_CELL_12_3 VDD VSS BL3 BLB3 WL12 SRAM_6T_CELL
XSRAM_6T_CELL_12_4 VDD VSS BL4 BLB4 WL12 SRAM_6T_CELL
XSRAM_6T_CELL_12_5 VDD VSS BL5 BLB5 WL12 SRAM_6T_CELL
XSRAM_6T_CELL_12_6 VDD VSS BL6 BLB6 WL12 SRAM_6T_CELL
XSRAM_6T_CELL_12_7 VDD VSS BL7 BLB7 WL12 SRAM_6T_CELL
XSRAM_6T_CELL_13_0 VDD VSS BL0 BLB0 WL13 SRAM_6T_CELL
XSRAM_6T_CELL_13_1 VDD VSS BL1 BLB1 WL13 SRAM_6T_CELL
XSRAM_6T_CELL_13_2 VDD VSS BL2 BLB2 WL13 SRAM_6T_CELL
XSRAM_6T_CELL_13_3 VDD VSS BL3 BLB3 WL13 SRAM_6T_CELL
XSRAM_6T_CELL_13_4 VDD VSS BL4 BLB4 WL13 SRAM_6T_CELL
XSRAM_6T_CELL_13_5 VDD VSS BL5 BLB5 WL13 SRAM_6T_CELL
XSRAM_6T_CELL_13_6 VDD VSS BL6 BLB6 WL13 SRAM_6T_CELL
XSRAM_6T_CELL_13_7 VDD VSS BL7 BLB7 WL13 SRAM_6T_CELL
XSRAM_6T_CELL_14_0 VDD VSS BL0 BLB0 WL14 SRAM_6T_CELL
XSRAM_6T_CELL_14_1 VDD VSS BL1 BLB1 WL14 SRAM_6T_CELL
XSRAM_6T_CELL_14_2 VDD VSS BL2 BLB2 WL14 SRAM_6T_CELL
XSRAM_6T_CELL_14_3 VDD VSS BL3 BLB3 WL14 SRAM_6T_CELL
XSRAM_6T_CELL_14_4 VDD VSS BL4 BLB4 WL14 SRAM_6T_CELL
XSRAM_6T_CELL_14_5 VDD VSS BL5 BLB5 WL14 SRAM_6T_CELL
XSRAM_6T_CELL_14_6 VDD VSS BL6 BLB6 WL14 SRAM_6T_CELL
XSRAM_6T_CELL_14_7 VDD VSS BL7 BLB7 WL14 SRAM_6T_CELL
XSRAM_6T_CELL_15_0 VDD VSS BL0 BLB0 WL15 SRAM_6T_CELL
XSRAM_6T_CELL_15_1 VDD VSS BL1 BLB1 WL15 SRAM_6T_CELL
XSRAM_6T_CELL_15_2 VDD VSS BL2 BLB2 WL15 SRAM_6T_CELL
XSRAM_6T_CELL_15_3 VDD VSS BL3 BLB3 WL15 SRAM_6T_CELL
XSRAM_6T_CELL_15_4 VDD VSS BL4 BLB4 WL15 SRAM_6T_CELL
XSRAM_6T_CELL_15_5 VDD VSS BL5 BLB5 WL15 SRAM_6T_CELL
XSRAM_6T_CELL_15_6 VDD VSS BL6 BLB6 WL15 SRAM_6T_CELL
XSRAM_6T_CELL_15_7 VDD VSS BL7 BLB7 WL15 SRAM_6T_CELL
.ends SRAM_6T_CORE_16x8

.subckt sram_17x1_replica_column VDD VSS RBL RBLB WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 WL16
.subckt Replica_CELL VDD VSS RBL RBLB WL
MPGL RBL WL Q VSS NMOS_VTG l=5e-08 w=1.35e-07
MPGR RBLB WL VDD VSS NMOS_VTG l=5e-08 w=1.35e-07
MPDL Q VDD VSS VSS NMOS_VTG l=5e-08 w=9e-08
MPUL Q VDD VDD VDD PMOS_VTG l=5e-08 w=9e-08
MPDR VDD Q VSS VSS NMOS_VTG l=5e-08 w=9e-08
MPUR VDD Q VDD VDD PMOS_VTG l=5e-08 w=9e-08
.ends Replica_CELL
XReplica_CELL_0 VDD VSS RBL RBLB WL0 Replica_CELL
XReplica_CELL_1 VDD VSS RBL RBLB WL1 Replica_CELL
XReplica_CELL_2 VDD VSS RBL RBLB WL2 Replica_CELL
XReplica_CELL_3 VDD VSS RBL RBLB WL3 Replica_CELL
XReplica_CELL_4 VDD VSS RBL RBLB WL4 Replica_CELL
XReplica_CELL_5 VDD VSS RBL RBLB WL5 Replica_CELL
XReplica_CELL_6 VDD VSS RBL RBLB WL6 Replica_CELL
XReplica_CELL_7 VDD VSS RBL RBLB WL7 Replica_CELL
XReplica_CELL_8 VDD VSS RBL RBLB WL8 Replica_CELL
XReplica_CELL_9 VDD VSS RBL RBLB WL9 Replica_CELL
XReplica_CELL_10 VDD VSS RBL RBLB WL10 Replica_CELL
XReplica_CELL_11 VDD VSS RBL RBLB WL11 Replica_CELL
XReplica_CELL_12 VDD VSS RBL RBLB WL12 Replica_CELL
XReplica_CELL_13 VDD VSS RBL RBLB WL13 Replica_CELL
XReplica_CELL_14 VDD VSS RBL RBLB WL14 Replica_CELL
XReplica_CELL_15 VDD VSS RBL RBLB WL15 Replica_CELL
XReplica_CELL_16 VDD VSS RBL RBLB WL16 Replica_CELL
.ends sram_17x1_replica_column

.subckt AND2 VDD VSS A B Z
.subckt PNAND2 VDD VSS A B Z
Mpnand2_pmos1 Z A VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpnand2_pmos2 Z B VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpnand2_nmos1 Z B net1 VSS NMOS_VTG l=5e-08 w=1.8e-07
Mpnand2_nmos2 net1 A VSS VSS NMOS_VTG l=5e-08 w=1.8e-07
.ends PNAND2

.subckt PINV VDD VSS A Z
Mpinv_pmos Z A VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpinv_nmos Z A VSS VSS NMOS_VTG l=5e-08 w=9e-08
.ends PINV
XPNAND3 VDD VSS A B zb_int PNAND2
XPINV VDD VSS zb_int Z PINV
.ends AND2

.subckt TIME VDD VSS clk csb web clk_buf clk_bar cs_bar cs we_bar we gated_clk_bar gated_clk_buf wl_en A0 A1 A2 A3 A_dff0 A_dff1 A_dff2 A_dff3 rbl rbl_delay rbl_delay_bar s_en w_en PRE
.subckt ADDR_DFF VDD VSS CLK A0 A1 A2 A3 A_dff0 A_dff1 A_dff2 A_dff3
.subckt DFF VDD VSS D Q CLK
.subckt PINV1 VDD VSS A Z
Mpinv_pmos Z A VDD VDD PMOS_VTG l=5e-08 w=5e-07
Mpinv_nmos Z A VSS VSS NMOS_VTG l=5e-08 w=2.5e-07
.ends PINV1

.subckt TRANSMISSION_GATE VDD VSS IN OUT CTR_P CTR_N
Mtranspmos OUT CTR_P IN VDD PMOS_VTG l=5e-08 w=5e-07
Mtransnmos IN CTR_N OUT VSS NMOS_VTG l=5e-08 w=2.5e-07
.ends TRANSMISSION_GATE
Xinv1_clk VDD VSS CLK CLKB PINV1
Xinv2_D VDD VSS D D_b PINV1
Xtg1 VDD VSS D_b z1 CLK CLKB TRANSMISSION_GATE
Xinv3 VDD VSS z1 z2 PINV1
Xinv4 VDD VSS z2 z3 PINV1
Xtg2 VDD VSS z3 z1 CLKB CLK TRANSMISSION_GATE
Xinv5 VDD VSS z2 z4 PINV1
Xtg3 VDD VSS z4 z5 CLKB CLK TRANSMISSION_GATE
Xinv6 VDD VSS z5 Q PINV1
Xinv7 VDD VSS Q QB PINV1
Xtg4 VDD VSS QB z5 CLK CLKB TRANSMISSION_GATE
.ends DFF
Xdff_0 VDD VSS A0 A_dff0 CLK DFF
Xdff_1 VDD VSS A1 A_dff1 CLK DFF
Xdff_2 VDD VSS A2 A_dff2 CLK DFF
Xdff_3 VDD VSS A3 A_dff3 CLK DFF
.ends ADDR_DFF

.subckt pdrive VDD VSS A Z
.subckt PINV1 VDD VSS A Z
Mpinv_pmos Z A VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpinv_nmos Z A VSS VSS NMOS_VTG l=5e-08 w=9e-08
.ends PINV1

.subckt PINV2 VDD VSS A Z
Mpinv_pmos Z A VDD VDD PMOS_VTG l=5e-08 w=8.1e-07
Mpinv_nmos Z A VSS VSS NMOS_VTG l=5e-08 w=2.7e-07
.ends PINV2

.subckt PINV3 VDD VSS A Z
Mpinv_pmos Z A VDD VDD PMOS_VTG l=5e-08 w=1.08e-06
Mpinv_nmos Z A VSS VSS NMOS_VTG l=5e-08 w=3.6e-07
.ends PINV3

.subckt PINV4 VDD VSS A Z
Mpinv_pmos Z A VDD VDD PMOS_VTG l=5e-08 w=1.69e-06
Mpinv_nmos Z A VSS VSS NMOS_VTG l=5e-08 w=5.6e-07
.ends PINV4
Xbuf_inv1 VDD VSS A zb1_node PINV1
Xbuf_inv2 VDD VSS zb1_node zb2_node PINV2
Xbuf_inv3 VDD VSS zb2_node zb3_node PINV3
Xbuf_inv4 VDD VSS zb3_node Z PINV4
.ends pdrive

.subckt PINV VDD VSS A Z
Mpinv_pmos Z A VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpinv_nmos Z A VSS VSS NMOS_VTG l=5e-08 w=9e-08
.ends PINV

.subckt DFF_BUF VDD VSS D Q QB CLK
.subckt DFF VDD VSS D Q CLK
.subckt PINV1 VDD VSS A Z
Mpinv_pmos Z A VDD VDD PMOS_VTG l=5e-08 w=5e-07
Mpinv_nmos Z A VSS VSS NMOS_VTG l=5e-08 w=2.5e-07
.ends PINV1

.subckt TRANSMISSION_GATE VDD VSS IN OUT CTR_P CTR_N
Mtranspmos OUT CTR_P IN VDD PMOS_VTG l=5e-08 w=5e-07
Mtransnmos IN CTR_N OUT VSS NMOS_VTG l=5e-08 w=2.5e-07
.ends TRANSMISSION_GATE
Xinv1_clk VDD VSS CLK CLKB PINV1
Xinv2_D VDD VSS D D_b PINV1
Xtg1 VDD VSS D_b z1 CLK CLKB TRANSMISSION_GATE
Xinv3 VDD VSS z1 z2 PINV1
Xinv4 VDD VSS z2 z3 PINV1
Xtg2 VDD VSS z3 z1 CLKB CLK TRANSMISSION_GATE
Xinv5 VDD VSS z2 z4 PINV1
Xtg3 VDD VSS z4 z5 CLKB CLK TRANSMISSION_GATE
Xinv6 VDD VSS z5 Q PINV1
Xinv7 VDD VSS Q QB PINV1
Xtg4 VDD VSS QB z5 CLK CLKB TRANSMISSION_GATE
.ends DFF

.subckt PINV1 VDD VSS A Z
Mpinv_pmos Z A VDD VDD PMOS_VTG l=5e-08 w=5.4e-07
Mpinv_nmos Z A VSS VSS NMOS_VTG l=5e-08 w=1.8e-07
.ends PINV1

.subckt PINV2 VDD VSS A Z
Mpinv_pmos Z A VDD VDD PMOS_VTG l=5e-08 w=1.08e-06
Mpinv_nmos Z A VSS VSS NMOS_VTG l=5e-08 w=3.6e-07
.ends PINV2
Xdff VDD VSS D qint CLK DFF
Xinv1 VDD VSS qint QB PINV1
Xinv2 VDD VSS QB Q PINV2
.ends DFF_BUF

.subckt AND2 VDD VSS A B Z
.subckt PNAND2 VDD VSS A B Z
Mpnand2_pmos1 Z A VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpnand2_pmos2 Z B VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpnand2_nmos1 Z B net1 VSS NMOS_VTG l=5e-08 w=1.8e-07
Mpnand2_nmos2 net1 A VSS VSS NMOS_VTG l=5e-08 w=1.8e-07
.ends PNAND2

.subckt PINV VDD VSS A Z
Mpinv_pmos Z A VDD VDD PMOS_VTG l=5e-08 w=1.62e-06
Mpinv_nmos Z A VSS VSS NMOS_VTG l=5e-08 w=5.4e-07
.ends PINV
XPNAND3 VDD VSS A B zb_int PNAND2
XPINV VDD VSS zb_int Z PINV
.ends AND2

.subckt wl_pdrive VDD VSS A Z
.subckt PINV1 VDD VSS A Z
Mpinv_pmos Z A VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpinv_nmos Z A VSS VSS NMOS_VTG l=5e-08 w=9e-08
.ends PINV1

.subckt PINV2 VDD VSS A Z
Mpinv_pmos Z A VDD VDD PMOS_VTG l=5e-08 w=1.35e-06
Mpinv_nmos Z A VSS VSS NMOS_VTG l=5e-08 w=4.5e-07
.ends PINV2
Xbuf_inv1 VDD VSS A zb1_node PINV1
Xbuf_inv2 VDD VSS zb1_node Z PINV2
.ends wl_pdrive

.subckt delay_chain VDD VSS in out
.subckt PINV1 VDD VSS A Z
Mpinv_pmos Z A VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpinv_nmos Z A VSS VSS NMOS_VTG l=5e-08 w=9e-08
.ends PINV1
Xdinv0 VDD VSS in dout_1 PINV1
Xdload_0_0 VDD VSS dout_1 n_0_0 PINV1
Xdload_0_1 VDD VSS dout_1 n_0_1 PINV1
Xdload_0_2 VDD VSS dout_1 n_0_2 PINV1
Xdload_0_3 VDD VSS dout_1 n_0_3 PINV1
Xdinv1 VDD VSS dout_1 dout_2 PINV1
Xdload_1_0 VDD VSS dout_2 n_1_0 PINV1
Xdload_1_1 VDD VSS dout_2 n_1_1 PINV1
Xdload_1_2 VDD VSS dout_2 n_1_2 PINV1
Xdload_1_3 VDD VSS dout_2 n_1_3 PINV1
Xdinv2 VDD VSS dout_2 dout_3 PINV1
Xdload_2_0 VDD VSS dout_3 n_2_0 PINV1
Xdload_2_1 VDD VSS dout_3 n_2_1 PINV1
Xdload_2_2 VDD VSS dout_3 n_2_2 PINV1
Xdload_2_3 VDD VSS dout_3 n_2_3 PINV1
Xdinv3 VDD VSS dout_3 dout_4 PINV1
Xdload_3_0 VDD VSS dout_4 n_3_0 PINV1
Xdload_3_1 VDD VSS dout_4 n_3_1 PINV1
Xdload_3_2 VDD VSS dout_4 n_3_2 PINV1
Xdload_3_3 VDD VSS dout_4 n_3_3 PINV1
Xdinv4 VDD VSS dout_4 dout_5 PINV1
Xdload_4_0 VDD VSS dout_5 n_4_0 PINV1
Xdload_4_1 VDD VSS dout_5 n_4_1 PINV1
Xdload_4_2 VDD VSS dout_5 n_4_2 PINV1
Xdload_4_3 VDD VSS dout_5 n_4_3 PINV1
Xdinv5 VDD VSS dout_5 dout_6 PINV1
Xdload_5_0 VDD VSS dout_6 n_5_0 PINV1
Xdload_5_1 VDD VSS dout_6 n_5_1 PINV1
Xdload_5_2 VDD VSS dout_6 n_5_2 PINV1
Xdload_5_3 VDD VSS dout_6 n_5_3 PINV1
Xdinv6 VDD VSS dout_6 dout_7 PINV1
Xdload_6_0 VDD VSS dout_7 n_6_0 PINV1
Xdload_6_1 VDD VSS dout_7 n_6_1 PINV1
Xdload_6_2 VDD VSS dout_7 n_6_2 PINV1
Xdload_6_3 VDD VSS dout_7 n_6_3 PINV1
Xdinv7 VDD VSS dout_7 dout_8 PINV1
Xdload_7_0 VDD VSS dout_8 n_7_0 PINV1
Xdload_7_1 VDD VSS dout_8 n_7_1 PINV1
Xdload_7_2 VDD VSS dout_8 n_7_2 PINV1
Xdload_7_3 VDD VSS dout_8 n_7_3 PINV1
Xdinv8 VDD VSS dout_8 out PINV1
Xdload_8_0 VDD VSS out n_8_0 PINV1
Xdload_8_1 VDD VSS out n_8_1 PINV1
Xdload_8_2 VDD VSS out n_8_2 PINV1
Xdload_8_3 VDD VSS out n_8_3 PINV1
.ends delay_chain

.subckt AND3 VDD VSS A B C Z
.subckt PNAND3 VDD VSS A B C Z
Mpnand3_pmos1 Z A VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpnand3_pmos2 Z B VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpnand3_pmos3 Z C VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpnand3_nmos1 Z A net1 VSS NMOS_VTG l=5e-08 w=1.8e-07
Mpnand3_nmos2 net1 B net2 VSS NMOS_VTG l=5e-08 w=1.8e-07
Mpnand3_nmos3 net2 C VSS VSS NMOS_VTG l=5e-08 w=1.8e-07
.ends PNAND3

.subckt PINV VDD VSS A Z
Mpinv_pmos Z A VDD VDD PMOS_VTG l=5e-08 w=1.08e-06
Mpinv_nmos Z A VSS VSS NMOS_VTG l=5e-08 w=3.6e-07
.ends PINV
XPNAND3 VDD VSS A B C zb_int PNAND3
XPINV VDD VSS zb_int Z PINV
.ends AND3

.subckt PNAND2 VDD VSS A B Z
Mpnand2_pmos1 Z A VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpnand2_pmos2 Z B VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpnand2_nmos1 Z B net1 VSS NMOS_VTG l=5e-08 w=1.8e-07
Mpnand2_nmos2 net1 A VSS VSS NMOS_VTG l=5e-08 w=1.8e-07
.ends PNAND2

.subckt pdrive2_for_pre VDD VSS A Z
.subckt PINV1 VDD VSS A Z
Mpinv_pmos Z A VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpinv_nmos Z A VSS VSS NMOS_VTG l=5e-08 w=9e-08
.ends PINV1

.subckt PINV2 VDD VSS A Z
Mpinv_pmos Z A VDD VDD PMOS_VTG l=5e-08 w=8.1e-07
Mpinv_nmos Z A VSS VSS NMOS_VTG l=5e-08 w=2.7e-07
.ends PINV2
Xbuf_inv1 VDD VSS A zb1_node PINV1
Xbuf_inv2 VDD VSS zb1_node Z PINV2
.ends pdrive2_for_pre
Xdff_buf_addr VDD VSS clk_buf A0 A1 A2 A3 A_dff0 A_dff1 A_dff2 A_dff3 ADDR_DFF
Xclkbuf VDD VSS clk clk_buf pdrive
Xinv_clk_bar VDD VSS clk_buf clk_bar PINV
Xdff_buf VDD VSS csb cs_bar cs clk_buf DFF_BUF
Xdff_buf1 VDD VSS web we_bar we clk_buf DFF_BUF
Xand2_gated_clk_bar VDD VSS cs clk_bar gated_clk_bar AND2
Xand2_gated_clk_buf VDD VSS cs clk_buf gated_clk_buf AND2
Xwl_en VDD VSS gated_clk_bar wl_en wl_pdrive
Xdelaychain VDD VSS rbl rbl_delay delay_chain
Xinv_rbl_delay_bar VDD VSS rbl_delay rbl_delay_bar PINV
Xw_en VDD VSS rbl_delay_bar gated_clk_bar we w_en AND3
Xs_en VDD VSS rbl_delay gated_clk_bar we_bar s_en AND3
Xpre_unbuf VDD VSS gated_clk_buf rbl_delay PRE_UNBUF PNAND2
Xpre VDD VSS PRE_UNBUF PRE pdrive2_for_pre
.ends TIME

.subckt DECODER_CASCADE VDD VSS A0 A1 A2 A3 WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15
.subckt DECODER3_8 VDD VSS EN A0 A1 A2 WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7
.subckt PINV VDD VSS A Z
Mpinv_pmos Z A VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpinv_nmos Z A VSS VSS NMOS_VTG l=5e-08 w=9e-08
.ends PINV

.subckt AND3 VDD VSS A B C Z
.subckt PNAND3 VDD VSS A B C Z
Mpnand3_pmos1 Z A VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpnand3_pmos2 Z B VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpnand3_pmos3 Z C VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpnand3_nmos1 Z A net1 VSS NMOS_VTG l=5e-08 w=1.8e-07
Mpnand3_nmos2 net1 B net2 VSS NMOS_VTG l=5e-08 w=1.8e-07
Mpnand3_nmos3 net2 C VSS VSS NMOS_VTG l=5e-08 w=1.8e-07
.ends PNAND3

.subckt PINV VDD VSS A Z
Mpinv_pmos Z A VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpinv_nmos Z A VSS VSS NMOS_VTG l=5e-08 w=9e-08
.ends PINV
XPNAND3 VDD VSS A B C zb_int PNAND3
XPINV VDD VSS zb_int Z PINV
.ends AND3

.subckt AND2 VDD VSS A B Z
.subckt PNAND2 VDD VSS A B Z
Mpnand2_pmos1 Z A VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpnand2_pmos2 Z B VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpnand2_nmos1 Z B net1 VSS NMOS_VTG l=5e-08 w=1.8e-07
Mpnand2_nmos2 net1 A VSS VSS NMOS_VTG l=5e-08 w=1.8e-07
.ends PNAND2

.subckt PINV VDD VSS A Z
Mpinv_pmos Z A VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpinv_nmos Z A VSS VSS NMOS_VTG l=5e-08 w=9e-08
.ends PINV
XPNAND3 VDD VSS A B zb_int PNAND2
XPINV VDD VSS zb_int Z PINV
.ends AND2
XINV_A1 VDD VSS A0 A0b PINV
XINV_A2 VDD VSS A1 A1b PINV
XINV_A3 VDD VSS A2 A2b PINV
XAND0 VDD VSS A0b A1b A2b WL0_pre AND3
XAND_EN0 VDD VSS WL0_pre EN WL0 AND2
XAND1 VDD VSS A0b A1b A2 WL1_pre AND3
XAND_EN1 VDD VSS WL1_pre EN WL1 AND2
XAND2 VDD VSS A0b A1 A2b WL2_pre AND3
XAND_EN2 VDD VSS WL2_pre EN WL2 AND2
XAND3 VDD VSS A0b A1 A2 WL3_pre AND3
XAND_EN3 VDD VSS WL3_pre EN WL3 AND2
XAND4 VDD VSS A0 A1b A2b WL4_pre AND3
XAND_EN4 VDD VSS WL4_pre EN WL4 AND2
XAND5 VDD VSS A0 A1b A2 WL5_pre AND3
XAND_EN5 VDD VSS WL5_pre EN WL5 AND2
XAND6 VDD VSS A0 A1 A2b WL6_pre AND3
XAND_EN6 VDD VSS WL6_pre EN WL6 AND2
XAND7 VDD VSS A0 A1 A2 WL7_pre AND3
XAND_EN7 VDD VSS WL7_pre EN WL7 AND2
.ends DECODER3_8
XDEC_0_0 VDD VSS VDD VSS VSS A3 EN_0_0_0 EN_0_0_1 EN_0_0_2 EN_0_0_3 EN_0_0_4 EN_0_0_5 EN_0_0_6 EN_0_0_7 DECODER3_8
XDEC_1_0 VDD VSS EN_0_0_0 A2 A1 A0 WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 DECODER3_8
XDEC_1_1 VDD VSS EN_0_0_1 A2 A1 A0 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 DECODER3_8
.ends DECODER_CASCADE

.subckt WORDLINEDRIVER VDD VSS A B Z
.subckt PNAND2 VDD VSS A B Z
Mpnand2_pmos1 Z A VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpnand2_pmos2 Z B VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpnand2_nmos1 Z B net1 VSS NMOS_VTG l=5e-08 w=1.8e-07
Mpnand2_nmos2 net1 A VSS VSS NMOS_VTG l=5e-08 w=1.8e-07
.ends PNAND2

.subckt PINV VDD VSS A Z
Mpinv_pmos Z A VDD VDD PMOS_VTG l=5e-08 w=5.4e-07
Mpinv_nmos Z A VSS VSS NMOS_VTG l=5e-08 w=1.8e-07
.ends PINV
XPNAND2 VDD VSS A B zb_int PNAND2
XPINV VDD VSS zb_int Z PINV
.ends WORDLINEDRIVER

.subckt D_LATCH VDD VSS D EN Q QB
.subckt PNAND2 VDD VSS A B Z
Mpnand2_pmos1 Z A VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpnand2_pmos2 Z B VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpnand2_nmos1 Z B net1 VSS NMOS_VTG l=5e-08 w=1.8e-07
Mpnand2_nmos2 net1 A VSS VSS NMOS_VTG l=5e-08 w=1.8e-07
.ends PNAND2

.subckt PINV VDD VSS A Z
Mpinv_pmos Z A VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
Mpinv_nmos Z A VSS VSS NMOS_VTG l=5e-08 w=1.8e-07
.ends PINV
XINV1 VDD VSS D DB PINV
XNAND1 VDD VSS D EN INT1 PNAND2
XNAND2 VDD VSS DB EN INT2 PNAND2
XNAND3 VDD VSS INT1 QB Q PNAND2
XNAND4 VDD VSS INT2 Q QB PNAND2
.ends D_LATCH

.subckt PRECHARGE VDD ENB BL BLB
M1 BL ENB VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
M2 BLB ENB VDD VDD PMOS_VTG l=5e-08 w=2.7e-07
M3 BL ENB BLB VDD PMOS_VTG l=5e-08 w=2.7e-07
.ends PRECHARGE

.subckt SENSEAMP VDD VSS EN IN INB Q QB
M1 Q QB net1 VSS NMOS_VTG l=5e-08 w=2.7e-07
M2 Q QB VDD VDD PMOS_VTG l=5e-08 w=5.4e-07
M3 QB Q net1 VSS NMOS_VTG l=5e-08 w=2.7e-07
M4 QB Q VDD VDD PMOS_VTG l=5e-08 w=5.4e-07
M5 Q EN IN VDD PMOS_VTG l=5e-08 w=7.2e-07
M6 QB EN INB VDD PMOS_VTG l=5e-08 w=7.2e-07
M7 net1 EN VSS VSS NMOS_VTG l=5e-08 w=2.7e-07
.ends SENSEAMP
VVDD VDD VSS 1.0V
VVSS VSS 0 0V
XSRAM_6T_CORE_16x8 VDD VSS BL0 BL1 BL2 BL3 BL4 BL5 BL6 BL7 BLB0 BLB1 BLB2 BLB3 BLB4 BLB5 BLB6 BLB7 WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 SRAM_6T_CORE_16x8
Xsram_17x1_replica_column VDD VSS RBL RBLB RWL WL0 WL1 WL2 WL3 WL4 WL5 WL6 WL7 WL8 WL9 WL10 WL11 WL12 WL13 WL14 WL15 sram_17x1_replica_column
XRWL VDD VSS wl_en VDD RWL AND2
XTIME VDD VSS clk csb web clk_buf clk_bar cs_bar cs we_bar we gated_clk_bar gated_clk_buf wl_en A0 A1 A2 A3 A_dff0 A_dff1 A_dff2 A_dff3 rbl rbl_delay rbl_delay_bar s_en w_en PRE TIME
XDECODER VDD VSS A_dff0 A_dff1 A_dff2 A_dff3 DEC_WL0 DEC_WL1 DEC_WL2 DEC_WL3 DEC_WL4 DEC_WL5 DEC_WL6 DEC_WL7 DEC_WL8 DEC_WL9 DEC_WL10 DEC_WL11 DEC_WL12 DEC_WL13 DEC_WL14 DEC_WL15 DECODER_CASCADE
XWL_DRV_0 VDD VSS DEC_WL0 WL_EN WL0 WORDLINEDRIVER
XWL_DRV_1 VDD VSS DEC_WL1 WL_EN WL1 WORDLINEDRIVER
XWL_DRV_2 VDD VSS DEC_WL2 WL_EN WL2 WORDLINEDRIVER
XWL_DRV_3 VDD VSS DEC_WL3 WL_EN WL3 WORDLINEDRIVER
XWL_DRV_4 VDD VSS DEC_WL4 WL_EN WL4 WORDLINEDRIVER
XWL_DRV_5 VDD VSS DEC_WL5 WL_EN WL5 WORDLINEDRIVER
XWL_DRV_6 VDD VSS DEC_WL6 WL_EN WL6 WORDLINEDRIVER
XWL_DRV_7 VDD VSS DEC_WL7 WL_EN WL7 WORDLINEDRIVER
XWL_DRV_8 VDD VSS DEC_WL8 WL_EN WL8 WORDLINEDRIVER
XWL_DRV_9 VDD VSS DEC_WL9 WL_EN WL9 WORDLINEDRIVER
XWL_DRV_10 VDD VSS DEC_WL10 WL_EN WL10 WORDLINEDRIVER
XWL_DRV_11 VDD VSS DEC_WL11 WL_EN WL11 WORDLINEDRIVER
XWL_DRV_12 VDD VSS DEC_WL12 WL_EN WL12 WORDLINEDRIVER
XWL_DRV_13 VDD VSS DEC_WL13 WL_EN WL13 WORDLINEDRIVER
XWL_DRV_14 VDD VSS DEC_WL14 WL_EN WL14 WORDLINEDRIVER
XWL_DRV_15 VDD VSS DEC_WL15 WL_EN WL15 WORDLINEDRIVER
XD_LATCH VDD VSS SA_Q7 S_EN OUT OUT_B D_LATCH
XPRECHARGE_0 VDD PRE BL0 BLB0 PRECHARGE
XPRECHARGE_1 VDD PRE BL1 BLB1 PRECHARGE
XPRECHARGE_2 VDD PRE BL2 BLB2 PRECHARGE
XPRECHARGE_3 VDD PRE BL3 BLB3 PRECHARGE
XPRECHARGE_4 VDD PRE BL4 BLB4 PRECHARGE
XPRECHARGE_5 VDD PRE BL5 BLB5 PRECHARGE
XPRECHARGE_6 VDD PRE BL6 BLB6 PRECHARGE
XPRECHARGE_7 VDD PRE BL7 BLB7 PRECHARGE
XPRECHARGE_RBL VDD PRE RBL RBLB PRECHARGE
XSENSEAMP_0 VDD VSS s_en BL0 BLB0 SA_Q0 SA_QB0 SENSEAMP
XSENSEAMP_1 VDD VSS s_en BL1 BLB1 SA_Q1 SA_QB1 SENSEAMP
XSENSEAMP_2 VDD VSS s_en BL2 BLB2 SA_Q2 SA_QB2 SENSEAMP
XSENSEAMP_3 VDD VSS s_en BL3 BLB3 SA_Q3 SA_QB3 SENSEAMP
XSENSEAMP_4 VDD VSS s_en BL4 BLB4 SA_Q4 SA_QB4 SENSEAMP
XSENSEAMP_5 VDD VSS s_en BL5 BLB5 SA_Q5 SA_QB5 SENSEAMP
XSENSEAMP_6 VDD VSS s_en BL6 BLB6 SA_Q6 SA_QB6 SENSEAMP
XSENSEAMP_7 VDD VSS s_en BL7 BLB7 SA_Q7 SA_QB7 SENSEAMP
VADDR_0 A0 VSS DC 0V PULSE(0V 1.0V 0.5ns 0.05ns 0.05ns 1.0ns 5ns)
VADDR_1 A1 VSS DC 0V PULSE(0V 1.0V 0.5ns 0.05ns 0.05ns 1.0ns 5ns)
VADDR_2 A2 VSS DC 0V PULSE(0V 1.0V 0.5ns 0.05ns 0.05ns 1.0ns 5ns)
VADDR_3 A3 VSS DC 0V PULSE(0V 1.0V 0.5ns 0.05ns 0.05ns 1.0ns 5ns)
VCLK clk VSS DC 0V PULSE(0V 1.0V 1.0ns 0.05ns 0.05ns 2.5ns 5ns)
VCSB csb VSS DC 0V PULSE(0V 1.0V 0ns 0.05ns 0.05ns 0.5ns 5ns)
VWEB web VSS DC 0V PULSE(0V 1.0V 0.5ns 0.05ns 0.05ns 4.9ns 5ns)
.options TEMP = 27C
.options TNOM = 27C
.ic V(A_dff0)=0V V(A_dff1)=0V V(A_dff2)=0V V(A_dff3)=0V V(BL0)=0V V(BL1)=0V V(BL2)=0V V(BL3)=0V V(BL4)=0V V(BL5)=0V V(BL6)=0V V(BL7)=0V V(RBL)=0V V(SA_Q0)=0V V(SA_Q1)=0V V(SA_Q2)=0V V(SA_Q3)=0V V(SA_Q4)=0V V(SA_Q5)=0V V(SA_Q6)=0V V(SA_Q7)=0V V(SA_QB0)=1.0V V(SA_QB1)=1.0V V(SA_QB2)=1.0V V(SA_QB3)=1.0V V(SA_QB4)=1.0V V(SA_QB5)=1.0V V(SA_QB6)=1.0V V(SA_QB7)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_0_0:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_0_0:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_0_1:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_0_1:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_0_2:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_0_2:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_0_3:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_0_3:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_0_4:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_0_4:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_0_5:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_0_5:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_0_6:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_0_6:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_0_7:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_0_7:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_10_0:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_10_0:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_10_1:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_10_1:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_10_2:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_10_2:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_10_3:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_10_3:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_10_4:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_10_4:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_10_5:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_10_5:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_10_6:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_10_6:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_10_7:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_10_7:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_11_0:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_11_0:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_11_1:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_11_1:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_11_2:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_11_2:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_11_3:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_11_3:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_11_4:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_11_4:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_11_5:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_11_5:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_11_6:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_11_6:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_11_7:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_11_7:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_12_0:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_12_0:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_12_1:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_12_1:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_12_2:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_12_2:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_12_3:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_12_3:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_12_4:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_12_4:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_12_5:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_12_5:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_12_6:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_12_6:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_12_7:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_12_7:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_13_0:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_13_0:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_13_1:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_13_1:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_13_2:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_13_2:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_13_3:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_13_3:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_13_4:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_13_4:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_13_5:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_13_5:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_13_6:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_13_6:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_13_7:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_13_7:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_14_0:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_14_0:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_14_1:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_14_1:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_14_2:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_14_2:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_14_3:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_14_3:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_14_4:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_14_4:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_14_5:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_14_5:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_14_6:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_14_6:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_14_7:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_14_7:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_15_0:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_15_0:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_15_1:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_15_1:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_15_2:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_15_2:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_15_3:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_15_3:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_15_4:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_15_4:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_15_5:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_15_5:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_15_6:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_15_6:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_15_7:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_15_7:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_1_0:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_1_0:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_1_1:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_1_1:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_1_2:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_1_2:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_1_3:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_1_3:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_1_4:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_1_4:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_1_5:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_1_5:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_1_6:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_1_6:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_1_7:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_1_7:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_2_0:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_2_0:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_2_1:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_2_1:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_2_2:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_2_2:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_2_3:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_2_3:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_2_4:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_2_4:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_2_5:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_2_5:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_2_6:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_2_6:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_2_7:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_2_7:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_3_0:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_3_0:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_3_1:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_3_1:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_3_2:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_3_2:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_3_3:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_3_3:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_3_4:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_3_4:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_3_5:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_3_5:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_3_6:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_3_6:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_3_7:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_3_7:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_4_0:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_4_0:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_4_1:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_4_1:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_4_2:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_4_2:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_4_3:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_4_3:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_4_4:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_4_4:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_4_5:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_4_5:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_4_6:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_4_6:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_4_7:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_4_7:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_5_0:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_5_0:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_5_1:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_5_1:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_5_2:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_5_2:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_5_3:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_5_3:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_5_4:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_5_4:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_5_5:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_5_5:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_5_6:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_5_6:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_5_7:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_5_7:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_6_0:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_6_0:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_6_1:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_6_1:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_6_2:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_6_2:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_6_3:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_6_3:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_6_4:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_6_4:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_6_5:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_6_5:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_6_6:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_6_6:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_6_7:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_6_7:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_7_0:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_7_0:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_7_1:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_7_1:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_7_2:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_7_2:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_7_3:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_7_3:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_7_4:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_7_4:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_7_5:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_7_5:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_7_6:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_7_6:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_7_7:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_7_7:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_8_0:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_8_0:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_8_1:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_8_1:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_8_2:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_8_2:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_8_3:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_8_3:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_8_4:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_8_4:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_8_5:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_8_5:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_8_6:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_8_6:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_8_7:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_8_7:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_9_0:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_9_0:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_9_1:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_9_1:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_9_2:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_9_2:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_9_3:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_9_3:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_9_4:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_9_4:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_9_5:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_9_5:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_9_6:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_9_6:QB)=1.0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_9_7:Q)=0V V(XSRAM_6T_CORE_16x8:XSRAM_6T_CELL_9_7:QB)=1.0V V(cs_bar)=1.0V V(we)=1.0V
.meas TRAN TPRCH TRIG V(PRE)=0.5 FALL=1 TARG V(BL7)=0.9 RISE=1
.meas TRAN TDECODER TRIG V(A_dff0)=0.5 RISE=1 TARG V(DEC_WL15)=0.5 RISE=1
.meas TRAN TWLDRV TRIG V(wl_en)=0.5 RISE=1 TARG V(WL15)=0.5 RISE=1
.meas TRAN TWL WHEN V(WL15)=0.5 RISE=1 
.meas TRAN TBL WHEN V(BL7)='V(BLB7)-0.25' FALL=1
.meas TRAN TSWING PARAM='TBL-TWL'
.meas TRAN TSA TRIG V(s_en)=0.5 RISE=1 TARG V(SA_Q7)=0.01 FALL=1
.meas TRAN Ts_en TRIG V(S_EN)=0.01 RISE=2 TARG V(S_EN)=0.5 RISE=1
.meas TRAN PAVG AVG {V(VDD)*I(VVDD)} FROM=0.0 TO=1e-08
.meas TRAN PDYN AVG {V(VDD)*I(VVDD)} FROM=4e-09 TO=6.000000000000001e-09
.meas TRAN PSTC AVG {V(VDD)*I(VVDD)} FROM=6.000000000000001e-09 TO=1e-08
.end
